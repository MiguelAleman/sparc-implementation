module decoder_32(output reg [31:0] Y, input [4:0] S, input enable);
	always @ (S, enable)
		begin
			// DEBUG			
			// $display("%b", enable);	
			if(!enable)
				case(S)
				5'b00000: Y = 32'b11111111111111111111111111111110;
				5'b00001: Y = 32'b11111111111111111111111111111101;
				5'b00010: Y = 32'b11111111111111111111111111111011;
				5'b00011: Y = 32'b11111111111111111111111111110111;
				5'b00100: Y = 32'b11111111111111111111111111101111;
				5'b00101: Y = 32'b11111111111111111111111111011111;
				5'b00110: Y = 32'b11111111111111111111111110111111;
				5'b00111: Y = 32'b11111111111111111111111101111111;
				5'b01000: Y = 32'b11111111111111111111111011111111;
				5'b01001: Y = 32'b11111111111111111111110111111111;
				5'b01010: Y = 32'b11111111111111111111101111111111;
				5'b01011: Y = 32'b11111111111111111111011111111111;
				5'b01100: Y = 32'b11111111111111111110111111111111;
				5'b01101: Y = 32'b11111111111111111101111111111111;
				5'b01110: Y = 32'b11111111111111111011111111111111;
				5'b01111: Y = 32'b11111111111111110111111111111111;
				5'b10000: Y = 32'b11111111111111101111111111111111;
				5'b10001: Y = 32'b11111111111111011111111111111111;
				5'b10010: Y = 32'b11111111111110111111111111111111;
				5'b10011: Y = 32'b11111111111101111111111111111111;
				5'b10100: Y = 32'b11111111111011111111111111111111;
				5'b10101: Y = 32'b11111111110111111111111111111111;
				5'b10110: Y = 32'b11111111101111111111111111111111;
				5'b10111: Y = 32'b11111111011111111111111111111111;
				5'b11000: Y = 32'b11111110111111111111111111111111;
				5'b11001: Y = 32'b11111101111111111111111111111111;
				5'b11010: Y = 32'b11111011111111111111111111111111;
				5'b11011: Y = 32'b11110111111111111111111111111111;
				5'b11100: Y = 32'b11101111111111111111111111111111;
				5'b11101: Y = 32'b11011111111111111111111111111111;
				5'b11110: Y = 32'b10111111111111111111111111111111;
				5'b11111: Y = 32'b01111111111111111111111111111111;
				endcase
			else
				Y = 32'b11111111111111111111111111111111;
		end 
endmodule